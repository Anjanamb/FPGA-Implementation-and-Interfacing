module clk_200hz (
    input clk_50mhz,
    output reg clk_200hz
);

reg [25:0] counter = 0;

always @(posedge clk_50mhz) begin
    if (counter == 124999) begin
        counter <= 0;
        clk_200hz <= ~clk_200hz;
    end
    else begin
        counter <= counter + 1;
    end
end

endmodule
